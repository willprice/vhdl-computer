------------------------------------------------------------------------------
-- @file <Name of the file>
-- @brief <TO ADD>
-- @detais <TO ADD>
-------------------------------------------------------------------------------

-- import std_logic from the IEEE library. Should be done for ALL VHDL files.
library IEEE;
use IEEE.std_logic_1164.all;

-- Module Entity Declaration
entity <name of the module> is
   generic (
      -- module generics like port widths go here
   );
   port(
      -- port list goes here
   )
end entity <name of the module>;

-- Module Architecture
architecture arch_rtl of <name of the module> is

   -- Signal declarations go here

begin
   
   -- The guts of the module go here.

end architecture arch_rtl;
