------------------------------------------------------------------------------
-- @file <Name of the file>
-- @brief <TO ADD>
-- @details <TO ADD>
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;

entity <name of the module> is
   generic (
      -- module generics like port widths go here
   );
   port(
      -- port list goes here
   )
end entity <name of the module>;

architecture arch_rtl of <name of the module> is

   -- Signal declarations go here

begin
   
   -- The guts of the module go here.

end architecture arch_rtl;
