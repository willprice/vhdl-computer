--
-- This is the common package file.
-- All common types, constants etc go in here.
--

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

package common_types is

end package;
